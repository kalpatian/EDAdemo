library verilog;
use verilog.vl_types.all;
entity MUXK_tb is
end MUXK_tb;
