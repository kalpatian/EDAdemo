library verilog;
use verilog.vl_types.all;
entity select4_1_tb is
end select4_1_tb;
