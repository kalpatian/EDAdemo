library verilog;
use verilog.vl_types.all;
entity CNT10_Changed_tb is
end CNT10_Changed_tb;
