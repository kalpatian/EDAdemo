library verilog;
use verilog.vl_types.all;
entity ADDSUB16_tb is
end ADDSUB16_tb;
