library verilog;
use verilog.vl_types.all;
entity tri_tb is
end tri_tb;
