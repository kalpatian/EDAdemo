library verilog;
use verilog.vl_types.all;
entity LS160_tb is
end LS160_tb;
