library verilog;
use verilog.vl_types.all;
entity CNT10_tb is
end CNT10_tb;
